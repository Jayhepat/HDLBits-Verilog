Build an XOR gate three ways, using an assign statement, a combinational always block, 
and a clocked always block. Note that the clocked always block produces a different circuit from the other two: There is a flip-flop so the output is delayed.

  CKT MODEL BLOCK: https://hdlbits.01xz.net/mw/images/4/40/Alwaysff.png
-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------

module top_module(
    input clk,
    input a,
    input b,
    output wire out_assign,
    output reg out_always_comb,
    output reg out_always_ff   );

endmodule
