Implement the following Circuit
CIRCUIT: https://hdlbits.01xz.net/wiki/File:Exams_m2014q4i.png

----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
module top_module(
  output out
);
  
  assign out = 1'b0;
  
  end module
