module top_module( input in, output out );
    
    assign out = !in;  // bitwise-NOT (~) and logical-NOT (!) operators, like C
endmodule
